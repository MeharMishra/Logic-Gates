// Code your design here
module nandgate(input a, input b, output c);
  assign c = ~(a & b);
endmodule