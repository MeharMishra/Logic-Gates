// Code your design here
module xorgate(input a, input b, output c);
  assign c = a ^ b;
endmodule