// Code your design here
module orgate(input a, input b, output c);
  assign c = a | b;
endmodule