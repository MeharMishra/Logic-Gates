// Code your design here
module notgate(input a, output c);
  assign c = !a;
endmodule